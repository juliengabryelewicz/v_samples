module main

fn greet(msg string) {
	println(msg)
}

fn main() {
	greet("Hello, world!")
}
